module MorraCinese(
  input primo [1:0], secondo [1:0], inizia,
  output manche [1:0], partita[1:0]
  );
   

endmodule
